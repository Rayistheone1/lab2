----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/25/2025 03:52:34 PM
-- Design Name: 
-- Module Name: sevenseg_decoder - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sevenseg_decoder is
    Port ( i_Hex : in STD_LOGIC_VECTOR (3 downto 0);
           o_seg_n : out STD_LOGIC_VECTOR (6 downto 0));
end sevenseg_decoder;

architecture Behavioral of sevenseg_decoder is
    signal w_sel: std_logic_vector (3 downto 0);

begin

w_sel(0) <= i_Hex(0);
w_sel(1) <= i_Hex(1);
w_sel(2) <= i_Hex(2);
w_sel(3) <= i_Hex(3);

with w_sel select
    o_seg_n <= "1000000" when "0000",
--        "1001111" when "0001",
        "1111001" when "0001", --flipped left/right
--        "0010010" when "0010", 
        "0100100" when "0010", --inverted all the bits
--        "0000110" when "0011", 
        "0110000" when "0011", --inverted and flipped all the bits
        "0011001" when "0100",
        "0010010" when "0101",
        "0000010" when "0110",
        "1111000" when "0111",
        "0000000" when "1000",
        "0011000" when "1001",
        "0001000" when "1010",
        "0000011" when "1011",
        "0100111" when "1100",
        "0100001" when "1101",
        "0000110" when "1110",
        "0001110" when "1111",
        "0000000" when others;


end Behavioral;
